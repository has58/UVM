// Simple Hello World module
module dut(dut_if dif);
endmodule


//---------------------------------------
// Interface Hello World
//---------------------------------------
interface dut_if(

);
endinterface
