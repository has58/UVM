// Simple adder/subtractor module
module dut(dut_if dif);
endmodule


//---------------------------------------
// Interface for the adder/subtractor DUT
//---------------------------------------
interface dut_if(

);
endinterface
